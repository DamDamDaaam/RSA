`timescale 1ns / 100ps

module Euclid(

);



endmodule
