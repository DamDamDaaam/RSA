`timescale 1ns / 100ps

module DecrypterOut (
    input wire clk,
    input wire rst
    );
    
    
    
endmodule
